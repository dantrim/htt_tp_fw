// SpyProtocol verilog include file.

// I chose these pretty arbitrarily. We can adjust as needed or add more
// valid metadata words.
parameter START_EVENT = 4'b1010;
parameter END_EVENT = 4'b0101;
